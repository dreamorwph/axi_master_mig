module a ();

sda
