module a ();

sd\
w23
